// Generator : SpinalHDL v1.10.1    git head : 2527c7c6b0fb0f95e5e1a5722a0be732b364ce43
// Component : SystolicArray2D
// Git hash  : cf1cfaa47c74a9bd373ec31b94c3beb4a5766bb1

`timescale 1ns/1ps 
module SystolicArray2D (
  input  wire          io_in_MatA_Bus_valid,
  output wire          io_in_MatA_Bus_ready,
  input  wire          io_in_MatA_Bus_payload_0_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_0_payload,
  input  wire          io_in_MatA_Bus_payload_1_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_1_payload,
  input  wire          io_in_MatA_Bus_payload_2_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_2_payload,
  input  wire          io_in_MatA_Bus_payload_3_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_3_payload,
  input  wire          io_in_MatA_Bus_payload_4_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_4_payload,
  input  wire          io_in_MatA_Bus_payload_5_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_5_payload,
  input  wire          io_in_MatA_Bus_payload_6_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_6_payload,
  input  wire          io_in_MatA_Bus_payload_7_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_7_payload,
  input  wire          io_in_MatA_Bus_payload_8_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_8_payload,
  input  wire          io_in_MatA_Bus_payload_9_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_9_payload,
  input  wire          io_in_MatA_Bus_payload_10_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_10_payload,
  input  wire          io_in_MatA_Bus_payload_11_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_11_payload,
  input  wire          io_in_MatA_Bus_payload_12_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_12_payload,
  input  wire          io_in_MatA_Bus_payload_13_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_13_payload,
  input  wire          io_in_MatA_Bus_payload_14_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_14_payload,
  input  wire          io_in_MatA_Bus_payload_15_valid,
  input  wire [15:0]   io_in_MatA_Bus_payload_15_payload,
  input  wire          io_in_MatB_Bus_valid,
  output wire          io_in_MatB_Bus_ready,
  input  wire          io_in_MatB_Bus_payload_0_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_0_payload,
  input  wire          io_in_MatB_Bus_payload_1_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_1_payload,
  input  wire          io_in_MatB_Bus_payload_2_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_2_payload,
  input  wire          io_in_MatB_Bus_payload_3_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_3_payload,
  input  wire          io_in_MatB_Bus_payload_4_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_4_payload,
  input  wire          io_in_MatB_Bus_payload_5_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_5_payload,
  input  wire          io_in_MatB_Bus_payload_6_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_6_payload,
  input  wire          io_in_MatB_Bus_payload_7_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_7_payload,
  input  wire          io_in_MatB_Bus_payload_8_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_8_payload,
  input  wire          io_in_MatB_Bus_payload_9_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_9_payload,
  input  wire          io_in_MatB_Bus_payload_10_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_10_payload,
  input  wire          io_in_MatB_Bus_payload_11_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_11_payload,
  input  wire          io_in_MatB_Bus_payload_12_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_12_payload,
  input  wire          io_in_MatB_Bus_payload_13_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_13_payload,
  input  wire          io_in_MatB_Bus_payload_14_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_14_payload,
  input  wire          io_in_MatB_Bus_payload_15_valid,
  input  wire [15:0]   io_in_MatB_Bus_payload_15_payload
);


  assign io_in_MatA_Bus_ready = 1'b1;
  assign io_in_MatB_Bus_ready = 1'b1;

endmodule
