// Generator : SpinalHDL v1.10.1    git head : 2527c7c6b0fb0f95e5e1a5722a0be732b364ce43
// Component : SystolicArray2D
// Git hash  : d927a680082e85a7bce9084e90db181aced08c49

`timescale 1ns/1ps 
module SystolicArray2D (
  input  wire          io_in_Mats_valid,
  output wire          io_in_Mats_ready,
  input  wire [15:0]   io_in_Mats_payload_A_0_data,
  input  wire          io_in_Mats_payload_A_0_Final,
  input  wire [15:0]   io_in_Mats_payload_A_1_data,
  input  wire          io_in_Mats_payload_A_1_Final,
  input  wire [15:0]   io_in_Mats_payload_A_2_data,
  input  wire          io_in_Mats_payload_A_2_Final,
  input  wire [15:0]   io_in_Mats_payload_B_0_data,
  input  wire          io_in_Mats_payload_B_0_Final,
  input  wire [15:0]   io_in_Mats_payload_B_1_data,
  input  wire          io_in_Mats_payload_B_1_Final,
  input  wire [15:0]   io_in_Mats_payload_B_2_data,
  input  wire          io_in_Mats_payload_B_2_Final,
  input  wire [15:0]   io_in_Mats_payload_B_3_data,
  input  wire          io_in_Mats_payload_B_3_Final,
  input  wire [15:0]   io_in_Mats_payload_B_4_data,
  input  wire          io_in_Mats_payload_B_4_Final,
  output wire          io_out_MatZ_valid,
  input  wire          io_out_MatZ_ready,
  output wire [31:0]   io_out_MatZ_payload_0_0,
  output wire [31:0]   io_out_MatZ_payload_0_1,
  output wire [31:0]   io_out_MatZ_payload_0_2,
  output wire [31:0]   io_out_MatZ_payload_0_3,
  output wire [31:0]   io_out_MatZ_payload_0_4,
  output wire [31:0]   io_out_MatZ_payload_1_0,
  output wire [31:0]   io_out_MatZ_payload_1_1,
  output wire [31:0]   io_out_MatZ_payload_1_2,
  output wire [31:0]   io_out_MatZ_payload_1_3,
  output wire [31:0]   io_out_MatZ_payload_1_4,
  output wire [31:0]   io_out_MatZ_payload_2_0,
  output wire [31:0]   io_out_MatZ_payload_2_1,
  output wire [31:0]   io_out_MatZ_payload_2_2,
  output wire [31:0]   io_out_MatZ_payload_2_3,
  output wire [31:0]   io_out_MatZ_payload_2_4,
  input  wire          clk,
  input  wire          resetn
);

  wire       [15:0]   systolicArray2DUnit_15_io_outA;
  wire                systolicArray2DUnit_15_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_15_io_outB;
  wire                systolicArray2DUnit_15_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_15_io_outZ;
  wire       [15:0]   systolicArray2DUnit_16_io_outA;
  wire                systolicArray2DUnit_16_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_16_io_outB;
  wire                systolicArray2DUnit_16_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_16_io_outZ;
  wire       [15:0]   systolicArray2DUnit_17_io_outA;
  wire                systolicArray2DUnit_17_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_17_io_outB;
  wire                systolicArray2DUnit_17_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_17_io_outZ;
  wire       [15:0]   systolicArray2DUnit_18_io_outA;
  wire                systolicArray2DUnit_18_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_18_io_outB;
  wire                systolicArray2DUnit_18_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_18_io_outZ;
  wire       [15:0]   systolicArray2DUnit_19_io_outA;
  wire                systolicArray2DUnit_19_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_19_io_outB;
  wire                systolicArray2DUnit_19_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_19_io_outZ;
  wire       [15:0]   systolicArray2DUnit_20_io_outA;
  wire                systolicArray2DUnit_20_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_20_io_outB;
  wire                systolicArray2DUnit_20_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_20_io_outZ;
  wire       [15:0]   systolicArray2DUnit_21_io_outA;
  wire                systolicArray2DUnit_21_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_21_io_outB;
  wire                systolicArray2DUnit_21_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_21_io_outZ;
  wire       [15:0]   systolicArray2DUnit_22_io_outA;
  wire                systolicArray2DUnit_22_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_22_io_outB;
  wire                systolicArray2DUnit_22_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_22_io_outZ;
  wire       [15:0]   systolicArray2DUnit_23_io_outA;
  wire                systolicArray2DUnit_23_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_23_io_outB;
  wire                systolicArray2DUnit_23_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_23_io_outZ;
  wire       [15:0]   systolicArray2DUnit_24_io_outA;
  wire                systolicArray2DUnit_24_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_24_io_outB;
  wire                systolicArray2DUnit_24_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_24_io_outZ;
  wire       [15:0]   systolicArray2DUnit_25_io_outA;
  wire                systolicArray2DUnit_25_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_25_io_outB;
  wire                systolicArray2DUnit_25_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_25_io_outZ;
  wire       [15:0]   systolicArray2DUnit_26_io_outA;
  wire                systolicArray2DUnit_26_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_26_io_outB;
  wire                systolicArray2DUnit_26_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_26_io_outZ;
  wire       [15:0]   systolicArray2DUnit_27_io_outA;
  wire                systolicArray2DUnit_27_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_27_io_outB;
  wire                systolicArray2DUnit_27_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_27_io_outZ;
  wire       [15:0]   systolicArray2DUnit_28_io_outA;
  wire                systolicArray2DUnit_28_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_28_io_outB;
  wire                systolicArray2DUnit_28_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_28_io_outZ;
  wire       [15:0]   systolicArray2DUnit_29_io_outA;
  wire                systolicArray2DUnit_29_io_outA_Final;
  wire       [15:0]   systolicArray2DUnit_29_io_outB;
  wire                systolicArray2DUnit_29_io_outB_Final;
  wire       [31:0]   systolicArray2DUnit_29_io_outZ;
  wire       [1:0]    _zz_Unit2buffer_ptr_0;
  wire       [1:0]    _zz_Unit2buffer_ptr_0_1;
  reg        [31:0]   _zz_io_out_MatZ_payload_0_0;
  reg        [31:0]   _zz_io_out_MatZ_payload_0_1;
  reg        [31:0]   _zz_io_out_MatZ_payload_0_2;
  reg        [31:0]   _zz_io_out_MatZ_payload_0_3;
  reg        [31:0]   _zz_io_out_MatZ_payload_0_4;
  reg        [31:0]   _zz_io_out_MatZ_payload_1_0;
  reg        [31:0]   _zz_io_out_MatZ_payload_1_1;
  reg        [31:0]   _zz_io_out_MatZ_payload_1_2;
  reg        [31:0]   _zz_io_out_MatZ_payload_1_3;
  reg        [31:0]   _zz_io_out_MatZ_payload_1_4;
  reg        [31:0]   _zz_io_out_MatZ_payload_2_0;
  reg        [31:0]   _zz_io_out_MatZ_payload_2_1;
  reg        [31:0]   _zz_io_out_MatZ_payload_2_2;
  reg        [31:0]   _zz_io_out_MatZ_payload_2_3;
  reg        [31:0]   _zz_io_out_MatZ_payload_2_4;
  reg                 _zz_io_out_MatZ_valid;
  wire                Go;
  wire       [15:0]   in_MatA_AfterDelay_0_data;
  wire                in_MatA_AfterDelay_0_Final;
  wire       [15:0]   in_MatA_AfterDelay_1_data;
  wire                in_MatA_AfterDelay_1_Final;
  wire       [15:0]   in_MatA_AfterDelay_2_data;
  wire                in_MatA_AfterDelay_2_Final;
  reg        [15:0]   io_in_Mats_payload_A_1_delay_1_data;
  reg                 io_in_Mats_payload_A_1_delay_1_Final;
  reg        [15:0]   io_in_Mats_payload_A_2_delay_1_data;
  reg                 io_in_Mats_payload_A_2_delay_1_Final;
  reg        [15:0]   io_in_Mats_payload_A_2_delay_2_data;
  reg                 io_in_Mats_payload_A_2_delay_2_Final;
  wire       [15:0]   in_MatB_AfterDelay_0_data;
  wire                in_MatB_AfterDelay_0_Final;
  wire       [15:0]   in_MatB_AfterDelay_1_data;
  wire                in_MatB_AfterDelay_1_Final;
  wire       [15:0]   in_MatB_AfterDelay_2_data;
  wire                in_MatB_AfterDelay_2_Final;
  wire       [15:0]   in_MatB_AfterDelay_3_data;
  wire                in_MatB_AfterDelay_3_Final;
  wire       [15:0]   in_MatB_AfterDelay_4_data;
  wire                in_MatB_AfterDelay_4_Final;
  reg        [15:0]   io_in_Mats_payload_B_1_delay_1_data;
  reg                 io_in_Mats_payload_B_1_delay_1_Final;
  reg        [15:0]   io_in_Mats_payload_B_2_delay_1_data;
  reg                 io_in_Mats_payload_B_2_delay_1_Final;
  reg        [15:0]   io_in_Mats_payload_B_2_delay_2_data;
  reg                 io_in_Mats_payload_B_2_delay_2_Final;
  reg        [15:0]   io_in_Mats_payload_B_3_delay_1_data;
  reg                 io_in_Mats_payload_B_3_delay_1_Final;
  reg        [15:0]   io_in_Mats_payload_B_3_delay_2_data;
  reg                 io_in_Mats_payload_B_3_delay_2_Final;
  reg        [15:0]   io_in_Mats_payload_B_3_delay_3_data;
  reg                 io_in_Mats_payload_B_3_delay_3_Final;
  reg        [15:0]   io_in_Mats_payload_B_4_delay_1_data;
  reg                 io_in_Mats_payload_B_4_delay_1_Final;
  reg        [15:0]   io_in_Mats_payload_B_4_delay_2_data;
  reg                 io_in_Mats_payload_B_4_delay_2_Final;
  reg        [15:0]   io_in_Mats_payload_B_4_delay_3_data;
  reg                 io_in_Mats_payload_B_4_delay_3_Final;
  reg        [15:0]   io_in_Mats_payload_B_4_delay_4_data;
  reg                 io_in_Mats_payload_B_4_delay_4_Final;
  wire       [15:0]   interconnect_outA_with_inA_0_0_data;
  wire                interconnect_outA_with_inA_0_0_Final;
  wire       [15:0]   interconnect_outA_with_inA_0_1_data;
  wire                interconnect_outA_with_inA_0_1_Final;
  wire       [15:0]   interconnect_outA_with_inA_0_2_data;
  wire                interconnect_outA_with_inA_0_2_Final;
  wire       [15:0]   interconnect_outA_with_inA_0_3_data;
  wire                interconnect_outA_with_inA_0_3_Final;
  wire       [15:0]   interconnect_outA_with_inA_0_4_data;
  wire                interconnect_outA_with_inA_0_4_Final;
  wire       [15:0]   interconnect_outA_with_inA_1_0_data;
  wire                interconnect_outA_with_inA_1_0_Final;
  wire       [15:0]   interconnect_outA_with_inA_1_1_data;
  wire                interconnect_outA_with_inA_1_1_Final;
  wire       [15:0]   interconnect_outA_with_inA_1_2_data;
  wire                interconnect_outA_with_inA_1_2_Final;
  wire       [15:0]   interconnect_outA_with_inA_1_3_data;
  wire                interconnect_outA_with_inA_1_3_Final;
  wire       [15:0]   interconnect_outA_with_inA_1_4_data;
  wire                interconnect_outA_with_inA_1_4_Final;
  wire       [15:0]   interconnect_outA_with_inA_2_0_data;
  wire                interconnect_outA_with_inA_2_0_Final;
  wire       [15:0]   interconnect_outA_with_inA_2_1_data;
  wire                interconnect_outA_with_inA_2_1_Final;
  wire       [15:0]   interconnect_outA_with_inA_2_2_data;
  wire                interconnect_outA_with_inA_2_2_Final;
  wire       [15:0]   interconnect_outA_with_inA_2_3_data;
  wire                interconnect_outA_with_inA_2_3_Final;
  wire       [15:0]   interconnect_outA_with_inA_2_4_data;
  wire                interconnect_outA_with_inA_2_4_Final;
  wire       [15:0]   interconnect_outB_with_inB_0_0_data;
  wire                interconnect_outB_with_inB_0_0_Final;
  wire       [15:0]   interconnect_outB_with_inB_0_1_data;
  wire                interconnect_outB_with_inB_0_1_Final;
  wire       [15:0]   interconnect_outB_with_inB_0_2_data;
  wire                interconnect_outB_with_inB_0_2_Final;
  wire       [15:0]   interconnect_outB_with_inB_0_3_data;
  wire                interconnect_outB_with_inB_0_3_Final;
  wire       [15:0]   interconnect_outB_with_inB_0_4_data;
  wire                interconnect_outB_with_inB_0_4_Final;
  wire       [15:0]   interconnect_outB_with_inB_1_0_data;
  wire                interconnect_outB_with_inB_1_0_Final;
  wire       [15:0]   interconnect_outB_with_inB_1_1_data;
  wire                interconnect_outB_with_inB_1_1_Final;
  wire       [15:0]   interconnect_outB_with_inB_1_2_data;
  wire                interconnect_outB_with_inB_1_2_Final;
  wire       [15:0]   interconnect_outB_with_inB_1_3_data;
  wire                interconnect_outB_with_inB_1_3_Final;
  wire       [15:0]   interconnect_outB_with_inB_1_4_data;
  wire                interconnect_outB_with_inB_1_4_Final;
  wire       [15:0]   interconnect_outB_with_inB_2_0_data;
  wire                interconnect_outB_with_inB_2_0_Final;
  wire       [15:0]   interconnect_outB_with_inB_2_1_data;
  wire                interconnect_outB_with_inB_2_1_Final;
  wire       [15:0]   interconnect_outB_with_inB_2_2_data;
  wire                interconnect_outB_with_inB_2_2_Final;
  wire       [15:0]   interconnect_outB_with_inB_2_3_data;
  wire                interconnect_outB_with_inB_2_3_Final;
  wire       [15:0]   interconnect_outB_with_inB_2_4_data;
  wire                interconnect_outB_with_inB_2_4_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_0_0_data;
  wire                out_MatZ_Bundle_wire_0_0_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_0_1_data;
  wire                out_MatZ_Bundle_wire_0_1_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_0_2_data;
  wire                out_MatZ_Bundle_wire_0_2_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_0_3_data;
  wire                out_MatZ_Bundle_wire_0_3_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_0_4_data;
  wire                out_MatZ_Bundle_wire_0_4_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_1_0_data;
  wire                out_MatZ_Bundle_wire_1_0_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_1_1_data;
  wire                out_MatZ_Bundle_wire_1_1_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_1_2_data;
  wire                out_MatZ_Bundle_wire_1_2_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_1_3_data;
  wire                out_MatZ_Bundle_wire_1_3_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_1_4_data;
  wire                out_MatZ_Bundle_wire_1_4_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_2_0_data;
  wire                out_MatZ_Bundle_wire_2_0_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_2_1_data;
  wire                out_MatZ_Bundle_wire_2_1_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_2_2_data;
  wire                out_MatZ_Bundle_wire_2_2_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_2_3_data;
  wire                out_MatZ_Bundle_wire_2_3_Final;
  wire       [31:0]   out_MatZ_Bundle_wire_2_4_data;
  wire                out_MatZ_Bundle_wire_2_4_Final;
  reg        [31:0]   buffer_array_0_data_0_0;
  reg        [31:0]   buffer_array_0_data_0_1;
  reg        [31:0]   buffer_array_0_data_0_2;
  wire       [31:0]   buffer_array_0_data_0_3;
  wire       [31:0]   buffer_array_0_data_0_4;
  reg        [31:0]   buffer_array_0_data_1_0;
  reg        [31:0]   buffer_array_0_data_1_1;
  reg        [31:0]   buffer_array_0_data_1_2;
  wire       [31:0]   buffer_array_0_data_1_3;
  wire       [31:0]   buffer_array_0_data_1_4;
  reg        [31:0]   buffer_array_0_data_2_0;
  reg        [31:0]   buffer_array_0_data_2_1;
  reg        [31:0]   buffer_array_0_data_2_2;
  wire       [31:0]   buffer_array_0_data_2_3;
  wire       [31:0]   buffer_array_0_data_2_4;
  reg                 buffer_array_0_Occupied;
  reg                 buffer_array_0_Valid;
  reg        [31:0]   buffer_array_1_data_0_0;
  reg        [31:0]   buffer_array_1_data_0_1;
  reg        [31:0]   buffer_array_1_data_0_2;
  wire       [31:0]   buffer_array_1_data_0_3;
  wire       [31:0]   buffer_array_1_data_0_4;
  reg        [31:0]   buffer_array_1_data_1_0;
  reg        [31:0]   buffer_array_1_data_1_1;
  reg        [31:0]   buffer_array_1_data_1_2;
  wire       [31:0]   buffer_array_1_data_1_3;
  wire       [31:0]   buffer_array_1_data_1_4;
  reg        [31:0]   buffer_array_1_data_2_0;
  reg        [31:0]   buffer_array_1_data_2_1;
  reg        [31:0]   buffer_array_1_data_2_2;
  wire       [31:0]   buffer_array_1_data_2_3;
  wire       [31:0]   buffer_array_1_data_2_4;
  reg                 buffer_array_1_Occupied;
  reg                 buffer_array_1_Valid;
  reg        [31:0]   buffer_array_2_data_0_0;
  reg        [31:0]   buffer_array_2_data_0_1;
  reg        [31:0]   buffer_array_2_data_0_2;
  wire       [31:0]   buffer_array_2_data_0_3;
  wire       [31:0]   buffer_array_2_data_0_4;
  reg        [31:0]   buffer_array_2_data_1_0;
  reg        [31:0]   buffer_array_2_data_1_1;
  reg        [31:0]   buffer_array_2_data_1_2;
  wire       [31:0]   buffer_array_2_data_1_3;
  wire       [31:0]   buffer_array_2_data_1_4;
  reg        [31:0]   buffer_array_2_data_2_0;
  reg        [31:0]   buffer_array_2_data_2_1;
  reg        [31:0]   buffer_array_2_data_2_2;
  wire       [31:0]   buffer_array_2_data_2_3;
  wire       [31:0]   buffer_array_2_data_2_4;
  reg                 buffer_array_2_Occupied;
  reg                 buffer_array_2_Valid;
  reg        [1:0]    Unit2buffer_ptr_0;
  reg        [1:0]    Unit2buffer_ptr_1;
  reg        [1:0]    Unit2buffer_ptr_2;
  wire       [1:0]    buffer_array_output_ptr;
  wire       [3:0]    _zz_1;
  wire                _zz_2;
  wire                _zz_3;
  wire                _zz_4;
  wire       [3:0]    _zz_5;
  wire                _zz_6;
  wire                _zz_7;
  wire                _zz_8;
  wire       [3:0]    _zz_9;
  wire                _zz_10;
  wire                _zz_11;
  wire                _zz_12;

  assign _zz_Unit2buffer_ptr_0 = (Unit2buffer_ptr_0 + 2'b01);
  assign _zz_Unit2buffer_ptr_0_1 = (Unit2buffer_ptr_0 + 2'b01);
  SystolicArray2DUnit systolicArray2DUnit_15 (
    .io_inA        (in_MatA_AfterDelay_0_data[15:0]     ), //i
    .io_inA_Final  (in_MatA_AfterDelay_0_Final          ), //i
    .io_inB        (in_MatB_AfterDelay_0_data[15:0]     ), //i
    .io_inB_Final  (in_MatB_AfterDelay_0_Final          ), //i
    .io_Go         (Go                                  ), //i
    .io_outA       (systolicArray2DUnit_15_io_outA[15:0]), //o
    .io_outA_Final (systolicArray2DUnit_15_io_outA_Final), //o
    .io_outB       (systolicArray2DUnit_15_io_outB[15:0]), //o
    .io_outB_Final (systolicArray2DUnit_15_io_outB_Final), //o
    .io_outZ       (systolicArray2DUnit_15_io_outZ[31:0]), //o
    .clk           (clk                                 ), //i
    .resetn        (resetn                              )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_16 (
    .io_inA        (interconnect_outA_with_inA_0_0_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_0_0_Final     ), //i
    .io_inB        (in_MatB_AfterDelay_1_data[15:0]          ), //i
    .io_inB_Final  (in_MatB_AfterDelay_1_Final               ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_16_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_16_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_16_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_16_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_16_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_17 (
    .io_inA        (interconnect_outA_with_inA_0_1_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_0_1_Final     ), //i
    .io_inB        (in_MatB_AfterDelay_2_data[15:0]          ), //i
    .io_inB_Final  (in_MatB_AfterDelay_2_Final               ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_17_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_17_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_17_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_17_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_17_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_18 (
    .io_inA        (interconnect_outA_with_inA_0_2_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_0_2_Final     ), //i
    .io_inB        (in_MatB_AfterDelay_3_data[15:0]          ), //i
    .io_inB_Final  (in_MatB_AfterDelay_3_Final               ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_18_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_18_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_18_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_18_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_18_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_19 (
    .io_inA        (interconnect_outA_with_inA_0_3_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_0_3_Final     ), //i
    .io_inB        (in_MatB_AfterDelay_4_data[15:0]          ), //i
    .io_inB_Final  (in_MatB_AfterDelay_4_Final               ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_19_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_19_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_19_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_19_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_19_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_20 (
    .io_inA        (in_MatA_AfterDelay_1_data[15:0]          ), //i
    .io_inA_Final  (in_MatA_AfterDelay_1_Final               ), //i
    .io_inB        (interconnect_outB_with_inB_0_0_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_0_0_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_20_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_20_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_20_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_20_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_20_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_21 (
    .io_inA        (interconnect_outA_with_inA_1_0_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_1_0_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_0_1_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_0_1_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_21_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_21_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_21_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_21_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_21_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_22 (
    .io_inA        (interconnect_outA_with_inA_1_1_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_1_1_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_0_2_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_0_2_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_22_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_22_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_22_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_22_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_22_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_23 (
    .io_inA        (interconnect_outA_with_inA_1_2_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_1_2_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_0_3_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_0_3_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_23_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_23_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_23_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_23_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_23_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_24 (
    .io_inA        (interconnect_outA_with_inA_1_3_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_1_3_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_0_4_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_0_4_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_24_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_24_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_24_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_24_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_24_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_25 (
    .io_inA        (in_MatA_AfterDelay_2_data[15:0]          ), //i
    .io_inA_Final  (in_MatA_AfterDelay_2_Final               ), //i
    .io_inB        (interconnect_outB_with_inB_1_0_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_1_0_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_25_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_25_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_25_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_25_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_25_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_26 (
    .io_inA        (interconnect_outA_with_inA_2_0_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_2_0_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_1_1_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_1_1_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_26_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_26_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_26_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_26_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_26_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_27 (
    .io_inA        (interconnect_outA_with_inA_2_1_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_2_1_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_1_2_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_1_2_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_27_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_27_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_27_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_27_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_27_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_28 (
    .io_inA        (interconnect_outA_with_inA_2_2_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_2_2_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_1_3_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_1_3_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_28_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_28_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_28_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_28_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_28_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  SystolicArray2DUnit systolicArray2DUnit_29 (
    .io_inA        (interconnect_outA_with_inA_2_3_data[15:0]), //i
    .io_inA_Final  (interconnect_outA_with_inA_2_3_Final     ), //i
    .io_inB        (interconnect_outB_with_inB_1_4_data[15:0]), //i
    .io_inB_Final  (interconnect_outB_with_inB_1_4_Final     ), //i
    .io_Go         (Go                                       ), //i
    .io_outA       (systolicArray2DUnit_29_io_outA[15:0]     ), //o
    .io_outA_Final (systolicArray2DUnit_29_io_outA_Final     ), //o
    .io_outB       (systolicArray2DUnit_29_io_outB[15:0]     ), //o
    .io_outB_Final (systolicArray2DUnit_29_io_outB_Final     ), //o
    .io_outZ       (systolicArray2DUnit_29_io_outZ[31:0]     ), //o
    .clk           (clk                                      ), //i
    .resetn        (resetn                                   )  //i
  );
  always @(*) begin
    case(buffer_array_output_ptr)
      2'b00 : begin
        _zz_io_out_MatZ_payload_0_0 = buffer_array_0_data_0_0;
        _zz_io_out_MatZ_payload_0_1 = buffer_array_0_data_0_1;
        _zz_io_out_MatZ_payload_0_2 = buffer_array_0_data_0_2;
        _zz_io_out_MatZ_payload_0_3 = buffer_array_0_data_0_3;
        _zz_io_out_MatZ_payload_0_4 = buffer_array_0_data_0_4;
        _zz_io_out_MatZ_payload_1_0 = buffer_array_0_data_1_0;
        _zz_io_out_MatZ_payload_1_1 = buffer_array_0_data_1_1;
        _zz_io_out_MatZ_payload_1_2 = buffer_array_0_data_1_2;
        _zz_io_out_MatZ_payload_1_3 = buffer_array_0_data_1_3;
        _zz_io_out_MatZ_payload_1_4 = buffer_array_0_data_1_4;
        _zz_io_out_MatZ_payload_2_0 = buffer_array_0_data_2_0;
        _zz_io_out_MatZ_payload_2_1 = buffer_array_0_data_2_1;
        _zz_io_out_MatZ_payload_2_2 = buffer_array_0_data_2_2;
        _zz_io_out_MatZ_payload_2_3 = buffer_array_0_data_2_3;
        _zz_io_out_MatZ_payload_2_4 = buffer_array_0_data_2_4;
        _zz_io_out_MatZ_valid = buffer_array_0_Valid;
      end
      2'b01 : begin
        _zz_io_out_MatZ_payload_0_0 = buffer_array_1_data_0_0;
        _zz_io_out_MatZ_payload_0_1 = buffer_array_1_data_0_1;
        _zz_io_out_MatZ_payload_0_2 = buffer_array_1_data_0_2;
        _zz_io_out_MatZ_payload_0_3 = buffer_array_1_data_0_3;
        _zz_io_out_MatZ_payload_0_4 = buffer_array_1_data_0_4;
        _zz_io_out_MatZ_payload_1_0 = buffer_array_1_data_1_0;
        _zz_io_out_MatZ_payload_1_1 = buffer_array_1_data_1_1;
        _zz_io_out_MatZ_payload_1_2 = buffer_array_1_data_1_2;
        _zz_io_out_MatZ_payload_1_3 = buffer_array_1_data_1_3;
        _zz_io_out_MatZ_payload_1_4 = buffer_array_1_data_1_4;
        _zz_io_out_MatZ_payload_2_0 = buffer_array_1_data_2_0;
        _zz_io_out_MatZ_payload_2_1 = buffer_array_1_data_2_1;
        _zz_io_out_MatZ_payload_2_2 = buffer_array_1_data_2_2;
        _zz_io_out_MatZ_payload_2_3 = buffer_array_1_data_2_3;
        _zz_io_out_MatZ_payload_2_4 = buffer_array_1_data_2_4;
        _zz_io_out_MatZ_valid = buffer_array_1_Valid;
      end
      default : begin
        _zz_io_out_MatZ_payload_0_0 = buffer_array_2_data_0_0;
        _zz_io_out_MatZ_payload_0_1 = buffer_array_2_data_0_1;
        _zz_io_out_MatZ_payload_0_2 = buffer_array_2_data_0_2;
        _zz_io_out_MatZ_payload_0_3 = buffer_array_2_data_0_3;
        _zz_io_out_MatZ_payload_0_4 = buffer_array_2_data_0_4;
        _zz_io_out_MatZ_payload_1_0 = buffer_array_2_data_1_0;
        _zz_io_out_MatZ_payload_1_1 = buffer_array_2_data_1_1;
        _zz_io_out_MatZ_payload_1_2 = buffer_array_2_data_1_2;
        _zz_io_out_MatZ_payload_1_3 = buffer_array_2_data_1_3;
        _zz_io_out_MatZ_payload_1_4 = buffer_array_2_data_1_4;
        _zz_io_out_MatZ_payload_2_0 = buffer_array_2_data_2_0;
        _zz_io_out_MatZ_payload_2_1 = buffer_array_2_data_2_1;
        _zz_io_out_MatZ_payload_2_2 = buffer_array_2_data_2_2;
        _zz_io_out_MatZ_payload_2_3 = buffer_array_2_data_2_3;
        _zz_io_out_MatZ_payload_2_4 = buffer_array_2_data_2_4;
        _zz_io_out_MatZ_valid = buffer_array_2_Valid;
      end
    endcase
  end

  assign Go = (io_out_MatZ_ready && io_in_Mats_valid);
  assign in_MatA_AfterDelay_0_data = io_in_Mats_payload_A_0_data;
  assign in_MatA_AfterDelay_0_Final = io_in_Mats_payload_A_0_Final;
  assign in_MatA_AfterDelay_1_data = io_in_Mats_payload_A_1_delay_1_data;
  assign in_MatA_AfterDelay_1_Final = io_in_Mats_payload_A_1_delay_1_Final;
  assign in_MatA_AfterDelay_2_data = io_in_Mats_payload_A_2_delay_2_data;
  assign in_MatA_AfterDelay_2_Final = io_in_Mats_payload_A_2_delay_2_Final;
  assign in_MatB_AfterDelay_0_data = io_in_Mats_payload_B_0_data;
  assign in_MatB_AfterDelay_0_Final = io_in_Mats_payload_B_0_Final;
  assign in_MatB_AfterDelay_1_data = io_in_Mats_payload_B_1_delay_1_data;
  assign in_MatB_AfterDelay_1_Final = io_in_Mats_payload_B_1_delay_1_Final;
  assign in_MatB_AfterDelay_2_data = io_in_Mats_payload_B_2_delay_2_data;
  assign in_MatB_AfterDelay_2_Final = io_in_Mats_payload_B_2_delay_2_Final;
  assign in_MatB_AfterDelay_3_data = io_in_Mats_payload_B_3_delay_3_data;
  assign in_MatB_AfterDelay_3_Final = io_in_Mats_payload_B_3_delay_3_Final;
  assign in_MatB_AfterDelay_4_data = io_in_Mats_payload_B_4_delay_4_data;
  assign in_MatB_AfterDelay_4_Final = io_in_Mats_payload_B_4_delay_4_Final;
  assign interconnect_outA_with_inA_0_0_data = systolicArray2DUnit_15_io_outA;
  assign interconnect_outA_with_inA_0_0_Final = systolicArray2DUnit_15_io_outA_Final;
  assign interconnect_outB_with_inB_0_0_data = systolicArray2DUnit_15_io_outB;
  assign interconnect_outB_with_inB_0_0_Final = systolicArray2DUnit_15_io_outB_Final;
  assign out_MatZ_Bundle_wire_0_0_data = systolicArray2DUnit_15_io_outZ;
  assign out_MatZ_Bundle_wire_0_0_Final = (systolicArray2DUnit_15_io_outA_Final && systolicArray2DUnit_15_io_outB_Final);
  assign interconnect_outA_with_inA_0_1_data = systolicArray2DUnit_16_io_outA;
  assign interconnect_outA_with_inA_0_1_Final = systolicArray2DUnit_16_io_outA_Final;
  assign interconnect_outB_with_inB_0_1_data = systolicArray2DUnit_16_io_outB;
  assign interconnect_outB_with_inB_0_1_Final = systolicArray2DUnit_16_io_outB_Final;
  assign out_MatZ_Bundle_wire_0_1_data = systolicArray2DUnit_16_io_outZ;
  assign out_MatZ_Bundle_wire_0_1_Final = (systolicArray2DUnit_16_io_outA_Final && systolicArray2DUnit_16_io_outB_Final);
  assign interconnect_outA_with_inA_0_2_data = systolicArray2DUnit_17_io_outA;
  assign interconnect_outA_with_inA_0_2_Final = systolicArray2DUnit_17_io_outA_Final;
  assign interconnect_outB_with_inB_0_2_data = systolicArray2DUnit_17_io_outB;
  assign interconnect_outB_with_inB_0_2_Final = systolicArray2DUnit_17_io_outB_Final;
  assign out_MatZ_Bundle_wire_0_2_data = systolicArray2DUnit_17_io_outZ;
  assign out_MatZ_Bundle_wire_0_2_Final = (systolicArray2DUnit_17_io_outA_Final && systolicArray2DUnit_17_io_outB_Final);
  assign interconnect_outA_with_inA_0_3_data = systolicArray2DUnit_18_io_outA;
  assign interconnect_outA_with_inA_0_3_Final = systolicArray2DUnit_18_io_outA_Final;
  assign interconnect_outB_with_inB_0_3_data = systolicArray2DUnit_18_io_outB;
  assign interconnect_outB_with_inB_0_3_Final = systolicArray2DUnit_18_io_outB_Final;
  assign out_MatZ_Bundle_wire_0_3_data = systolicArray2DUnit_18_io_outZ;
  assign out_MatZ_Bundle_wire_0_3_Final = (systolicArray2DUnit_18_io_outA_Final && systolicArray2DUnit_18_io_outB_Final);
  assign interconnect_outA_with_inA_0_4_data = systolicArray2DUnit_19_io_outA;
  assign interconnect_outA_with_inA_0_4_Final = systolicArray2DUnit_19_io_outA_Final;
  assign interconnect_outB_with_inB_0_4_data = systolicArray2DUnit_19_io_outB;
  assign interconnect_outB_with_inB_0_4_Final = systolicArray2DUnit_19_io_outB_Final;
  assign out_MatZ_Bundle_wire_0_4_data = systolicArray2DUnit_19_io_outZ;
  assign out_MatZ_Bundle_wire_0_4_Final = (systolicArray2DUnit_19_io_outA_Final && systolicArray2DUnit_19_io_outB_Final);
  assign interconnect_outA_with_inA_1_0_data = systolicArray2DUnit_20_io_outA;
  assign interconnect_outA_with_inA_1_0_Final = systolicArray2DUnit_20_io_outA_Final;
  assign interconnect_outB_with_inB_1_0_data = systolicArray2DUnit_20_io_outB;
  assign interconnect_outB_with_inB_1_0_Final = systolicArray2DUnit_20_io_outB_Final;
  assign out_MatZ_Bundle_wire_1_0_data = systolicArray2DUnit_20_io_outZ;
  assign out_MatZ_Bundle_wire_1_0_Final = (systolicArray2DUnit_20_io_outA_Final && systolicArray2DUnit_20_io_outB_Final);
  assign interconnect_outA_with_inA_1_1_data = systolicArray2DUnit_21_io_outA;
  assign interconnect_outA_with_inA_1_1_Final = systolicArray2DUnit_21_io_outA_Final;
  assign interconnect_outB_with_inB_1_1_data = systolicArray2DUnit_21_io_outB;
  assign interconnect_outB_with_inB_1_1_Final = systolicArray2DUnit_21_io_outB_Final;
  assign out_MatZ_Bundle_wire_1_1_data = systolicArray2DUnit_21_io_outZ;
  assign out_MatZ_Bundle_wire_1_1_Final = (systolicArray2DUnit_21_io_outA_Final && systolicArray2DUnit_21_io_outB_Final);
  assign interconnect_outA_with_inA_1_2_data = systolicArray2DUnit_22_io_outA;
  assign interconnect_outA_with_inA_1_2_Final = systolicArray2DUnit_22_io_outA_Final;
  assign interconnect_outB_with_inB_1_2_data = systolicArray2DUnit_22_io_outB;
  assign interconnect_outB_with_inB_1_2_Final = systolicArray2DUnit_22_io_outB_Final;
  assign out_MatZ_Bundle_wire_1_2_data = systolicArray2DUnit_22_io_outZ;
  assign out_MatZ_Bundle_wire_1_2_Final = (systolicArray2DUnit_22_io_outA_Final && systolicArray2DUnit_22_io_outB_Final);
  assign interconnect_outA_with_inA_1_3_data = systolicArray2DUnit_23_io_outA;
  assign interconnect_outA_with_inA_1_3_Final = systolicArray2DUnit_23_io_outA_Final;
  assign interconnect_outB_with_inB_1_3_data = systolicArray2DUnit_23_io_outB;
  assign interconnect_outB_with_inB_1_3_Final = systolicArray2DUnit_23_io_outB_Final;
  assign out_MatZ_Bundle_wire_1_3_data = systolicArray2DUnit_23_io_outZ;
  assign out_MatZ_Bundle_wire_1_3_Final = (systolicArray2DUnit_23_io_outA_Final && systolicArray2DUnit_23_io_outB_Final);
  assign interconnect_outA_with_inA_1_4_data = systolicArray2DUnit_24_io_outA;
  assign interconnect_outA_with_inA_1_4_Final = systolicArray2DUnit_24_io_outA_Final;
  assign interconnect_outB_with_inB_1_4_data = systolicArray2DUnit_24_io_outB;
  assign interconnect_outB_with_inB_1_4_Final = systolicArray2DUnit_24_io_outB_Final;
  assign out_MatZ_Bundle_wire_1_4_data = systolicArray2DUnit_24_io_outZ;
  assign out_MatZ_Bundle_wire_1_4_Final = (systolicArray2DUnit_24_io_outA_Final && systolicArray2DUnit_24_io_outB_Final);
  assign interconnect_outA_with_inA_2_0_data = systolicArray2DUnit_25_io_outA;
  assign interconnect_outA_with_inA_2_0_Final = systolicArray2DUnit_25_io_outA_Final;
  assign interconnect_outB_with_inB_2_0_data = systolicArray2DUnit_25_io_outB;
  assign interconnect_outB_with_inB_2_0_Final = systolicArray2DUnit_25_io_outB_Final;
  assign out_MatZ_Bundle_wire_2_0_data = systolicArray2DUnit_25_io_outZ;
  assign out_MatZ_Bundle_wire_2_0_Final = (systolicArray2DUnit_25_io_outA_Final && systolicArray2DUnit_25_io_outB_Final);
  assign interconnect_outA_with_inA_2_1_data = systolicArray2DUnit_26_io_outA;
  assign interconnect_outA_with_inA_2_1_Final = systolicArray2DUnit_26_io_outA_Final;
  assign interconnect_outB_with_inB_2_1_data = systolicArray2DUnit_26_io_outB;
  assign interconnect_outB_with_inB_2_1_Final = systolicArray2DUnit_26_io_outB_Final;
  assign out_MatZ_Bundle_wire_2_1_data = systolicArray2DUnit_26_io_outZ;
  assign out_MatZ_Bundle_wire_2_1_Final = (systolicArray2DUnit_26_io_outA_Final && systolicArray2DUnit_26_io_outB_Final);
  assign interconnect_outA_with_inA_2_2_data = systolicArray2DUnit_27_io_outA;
  assign interconnect_outA_with_inA_2_2_Final = systolicArray2DUnit_27_io_outA_Final;
  assign interconnect_outB_with_inB_2_2_data = systolicArray2DUnit_27_io_outB;
  assign interconnect_outB_with_inB_2_2_Final = systolicArray2DUnit_27_io_outB_Final;
  assign out_MatZ_Bundle_wire_2_2_data = systolicArray2DUnit_27_io_outZ;
  assign out_MatZ_Bundle_wire_2_2_Final = (systolicArray2DUnit_27_io_outA_Final && systolicArray2DUnit_27_io_outB_Final);
  assign interconnect_outA_with_inA_2_3_data = systolicArray2DUnit_28_io_outA;
  assign interconnect_outA_with_inA_2_3_Final = systolicArray2DUnit_28_io_outA_Final;
  assign interconnect_outB_with_inB_2_3_data = systolicArray2DUnit_28_io_outB;
  assign interconnect_outB_with_inB_2_3_Final = systolicArray2DUnit_28_io_outB_Final;
  assign out_MatZ_Bundle_wire_2_3_data = systolicArray2DUnit_28_io_outZ;
  assign out_MatZ_Bundle_wire_2_3_Final = (systolicArray2DUnit_28_io_outA_Final && systolicArray2DUnit_28_io_outB_Final);
  assign interconnect_outA_with_inA_2_4_data = systolicArray2DUnit_29_io_outA;
  assign interconnect_outA_with_inA_2_4_Final = systolicArray2DUnit_29_io_outA_Final;
  assign interconnect_outB_with_inB_2_4_data = systolicArray2DUnit_29_io_outB;
  assign interconnect_outB_with_inB_2_4_Final = systolicArray2DUnit_29_io_outB_Final;
  assign out_MatZ_Bundle_wire_2_4_data = systolicArray2DUnit_29_io_outZ;
  assign out_MatZ_Bundle_wire_2_4_Final = (systolicArray2DUnit_29_io_outA_Final && systolicArray2DUnit_29_io_outB_Final);
  assign buffer_array_0_data_0_3 = 32'h00000000;
  assign buffer_array_0_data_0_4 = 32'h00000000;
  assign buffer_array_0_data_1_3 = 32'h00000000;
  assign buffer_array_0_data_1_4 = 32'h00000000;
  assign buffer_array_0_data_2_3 = 32'h00000000;
  assign buffer_array_0_data_2_4 = 32'h00000000;
  assign buffer_array_1_data_0_3 = 32'h00000000;
  assign buffer_array_1_data_0_4 = 32'h00000000;
  assign buffer_array_1_data_1_3 = 32'h00000000;
  assign buffer_array_1_data_1_4 = 32'h00000000;
  assign buffer_array_1_data_2_3 = 32'h00000000;
  assign buffer_array_1_data_2_4 = 32'h00000000;
  assign buffer_array_2_data_0_3 = 32'h00000000;
  assign buffer_array_2_data_0_4 = 32'h00000000;
  assign buffer_array_2_data_1_3 = 32'h00000000;
  assign buffer_array_2_data_1_4 = 32'h00000000;
  assign buffer_array_2_data_2_3 = 32'h00000000;
  assign buffer_array_2_data_2_4 = 32'h00000000;
  assign buffer_array_output_ptr = 2'b00;
  assign _zz_1 = ({3'd0,1'b1} <<< Unit2buffer_ptr_0);
  assign _zz_2 = _zz_1[0];
  assign _zz_3 = _zz_1[1];
  assign _zz_4 = _zz_1[2];
  assign _zz_5 = ({3'd0,1'b1} <<< Unit2buffer_ptr_1);
  assign _zz_6 = _zz_5[0];
  assign _zz_7 = _zz_5[1];
  assign _zz_8 = _zz_5[2];
  assign _zz_9 = ({3'd0,1'b1} <<< Unit2buffer_ptr_2);
  assign _zz_10 = _zz_9[0];
  assign _zz_11 = _zz_9[1];
  assign _zz_12 = _zz_9[2];
  assign io_out_MatZ_payload_0_0 = _zz_io_out_MatZ_payload_0_0;
  assign io_out_MatZ_payload_0_1 = _zz_io_out_MatZ_payload_0_1;
  assign io_out_MatZ_payload_0_2 = _zz_io_out_MatZ_payload_0_2;
  assign io_out_MatZ_payload_0_3 = _zz_io_out_MatZ_payload_0_3;
  assign io_out_MatZ_payload_0_4 = _zz_io_out_MatZ_payload_0_4;
  assign io_out_MatZ_payload_1_0 = _zz_io_out_MatZ_payload_1_0;
  assign io_out_MatZ_payload_1_1 = _zz_io_out_MatZ_payload_1_1;
  assign io_out_MatZ_payload_1_2 = _zz_io_out_MatZ_payload_1_2;
  assign io_out_MatZ_payload_1_3 = _zz_io_out_MatZ_payload_1_3;
  assign io_out_MatZ_payload_1_4 = _zz_io_out_MatZ_payload_1_4;
  assign io_out_MatZ_payload_2_0 = _zz_io_out_MatZ_payload_2_0;
  assign io_out_MatZ_payload_2_1 = _zz_io_out_MatZ_payload_2_1;
  assign io_out_MatZ_payload_2_2 = _zz_io_out_MatZ_payload_2_2;
  assign io_out_MatZ_payload_2_3 = _zz_io_out_MatZ_payload_2_3;
  assign io_out_MatZ_payload_2_4 = _zz_io_out_MatZ_payload_2_4;
  assign io_out_MatZ_valid = _zz_io_out_MatZ_valid;
  assign io_in_Mats_ready = io_out_MatZ_ready;
  always @(posedge clk) begin
    if(Go) begin
      io_in_Mats_payload_A_1_delay_1_data <= io_in_Mats_payload_A_1_data;
      io_in_Mats_payload_A_1_delay_1_Final <= io_in_Mats_payload_A_1_Final;
    end
    if(Go) begin
      io_in_Mats_payload_A_2_delay_1_data <= io_in_Mats_payload_A_2_data;
      io_in_Mats_payload_A_2_delay_1_Final <= io_in_Mats_payload_A_2_Final;
    end
    if(Go) begin
      io_in_Mats_payload_A_2_delay_2_data <= io_in_Mats_payload_A_2_delay_1_data;
      io_in_Mats_payload_A_2_delay_2_Final <= io_in_Mats_payload_A_2_delay_1_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_1_delay_1_data <= io_in_Mats_payload_B_1_data;
      io_in_Mats_payload_B_1_delay_1_Final <= io_in_Mats_payload_B_1_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_2_delay_1_data <= io_in_Mats_payload_B_2_data;
      io_in_Mats_payload_B_2_delay_1_Final <= io_in_Mats_payload_B_2_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_2_delay_2_data <= io_in_Mats_payload_B_2_delay_1_data;
      io_in_Mats_payload_B_2_delay_2_Final <= io_in_Mats_payload_B_2_delay_1_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_3_delay_1_data <= io_in_Mats_payload_B_3_data;
      io_in_Mats_payload_B_3_delay_1_Final <= io_in_Mats_payload_B_3_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_3_delay_2_data <= io_in_Mats_payload_B_3_delay_1_data;
      io_in_Mats_payload_B_3_delay_2_Final <= io_in_Mats_payload_B_3_delay_1_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_3_delay_3_data <= io_in_Mats_payload_B_3_delay_2_data;
      io_in_Mats_payload_B_3_delay_3_Final <= io_in_Mats_payload_B_3_delay_2_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_4_delay_1_data <= io_in_Mats_payload_B_4_data;
      io_in_Mats_payload_B_4_delay_1_Final <= io_in_Mats_payload_B_4_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_4_delay_2_data <= io_in_Mats_payload_B_4_delay_1_data;
      io_in_Mats_payload_B_4_delay_2_Final <= io_in_Mats_payload_B_4_delay_1_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_4_delay_3_data <= io_in_Mats_payload_B_4_delay_2_data;
      io_in_Mats_payload_B_4_delay_3_Final <= io_in_Mats_payload_B_4_delay_2_Final;
    end
    if(Go) begin
      io_in_Mats_payload_B_4_delay_4_data <= io_in_Mats_payload_B_4_delay_3_data;
      io_in_Mats_payload_B_4_delay_4_Final <= io_in_Mats_payload_B_4_delay_3_Final;
    end
  end

  always @(posedge clk or negedge resetn) begin
    if(!resetn) begin
      buffer_array_0_data_0_0 <= 32'h00000000;
      buffer_array_0_data_0_1 <= 32'h00000000;
      buffer_array_0_data_0_2 <= 32'h00000000;
      buffer_array_0_data_1_0 <= 32'h00000000;
      buffer_array_0_data_1_1 <= 32'h00000000;
      buffer_array_0_data_1_2 <= 32'h00000000;
      buffer_array_0_data_2_0 <= 32'h00000000;
      buffer_array_0_data_2_1 <= 32'h00000000;
      buffer_array_0_data_2_2 <= 32'h00000000;
      buffer_array_0_Occupied <= 1'b0;
      buffer_array_0_Valid <= 1'b0;
      buffer_array_1_data_0_0 <= 32'h00000000;
      buffer_array_1_data_0_1 <= 32'h00000000;
      buffer_array_1_data_0_2 <= 32'h00000000;
      buffer_array_1_data_1_0 <= 32'h00000000;
      buffer_array_1_data_1_1 <= 32'h00000000;
      buffer_array_1_data_1_2 <= 32'h00000000;
      buffer_array_1_data_2_0 <= 32'h00000000;
      buffer_array_1_data_2_1 <= 32'h00000000;
      buffer_array_1_data_2_2 <= 32'h00000000;
      buffer_array_1_Occupied <= 1'b0;
      buffer_array_1_Valid <= 1'b0;
      buffer_array_2_data_0_0 <= 32'h00000000;
      buffer_array_2_data_0_1 <= 32'h00000000;
      buffer_array_2_data_0_2 <= 32'h00000000;
      buffer_array_2_data_1_0 <= 32'h00000000;
      buffer_array_2_data_1_1 <= 32'h00000000;
      buffer_array_2_data_1_2 <= 32'h00000000;
      buffer_array_2_data_2_0 <= 32'h00000000;
      buffer_array_2_data_2_1 <= 32'h00000000;
      buffer_array_2_data_2_2 <= 32'h00000000;
      buffer_array_2_Occupied <= 1'b0;
      buffer_array_2_Valid <= 1'b0;
      Unit2buffer_ptr_0 <= 2'b00;
      Unit2buffer_ptr_1 <= 2'b00;
      Unit2buffer_ptr_2 <= 2'b00;
    end else begin
      if(Go) begin
        Unit2buffer_ptr_2 <= Unit2buffer_ptr_1;
        Unit2buffer_ptr_1 <= Unit2buffer_ptr_0;
        if(out_MatZ_Bundle_wire_0_0_Final) begin
          Unit2buffer_ptr_0 <= ((2'b11 <= _zz_Unit2buffer_ptr_0) ? _zz_Unit2buffer_ptr_0_1 : 2'b00);
          if(_zz_2) begin
            buffer_array_0_Occupied <= 1'b1;
          end
          if(_zz_3) begin
            buffer_array_1_Occupied <= 1'b1;
          end
          if(_zz_4) begin
            buffer_array_2_Occupied <= 1'b1;
          end
        end
        if(out_MatZ_Bundle_wire_2_4_Final) begin
          if(_zz_2) begin
            buffer_array_0_Valid <= 1'b1;
          end
          if(_zz_3) begin
            buffer_array_1_Valid <= 1'b1;
          end
          if(_zz_4) begin
            buffer_array_2_Valid <= 1'b1;
          end
        end else begin
          if(_zz_2) begin
            buffer_array_0_Valid <= 1'b0;
          end
          if(_zz_3) begin
            buffer_array_1_Valid <= 1'b0;
          end
          if(_zz_4) begin
            buffer_array_2_Valid <= 1'b0;
          end
        end
        if(buffer_array_0_Occupied) begin
          if(out_MatZ_Bundle_wire_0_0_Final) begin
            if(_zz_2) begin
              buffer_array_0_data_0_0 <= out_MatZ_Bundle_wire_0_0_data;
            end
            if(_zz_3) begin
              buffer_array_1_data_0_0 <= out_MatZ_Bundle_wire_0_0_data;
            end
            if(_zz_4) begin
              buffer_array_2_data_0_0 <= out_MatZ_Bundle_wire_0_0_data;
            end
          end
          if(buffer_array_0_Valid) begin
            buffer_array_0_Valid <= 1'b0;
            buffer_array_0_Occupied <= 1'b0;
          end
        end
        if(buffer_array_1_Occupied) begin
          if(out_MatZ_Bundle_wire_0_1_Final) begin
            if(_zz_6) begin
              buffer_array_0_data_0_1 <= out_MatZ_Bundle_wire_0_1_data;
            end
            if(_zz_7) begin
              buffer_array_1_data_0_1 <= out_MatZ_Bundle_wire_0_1_data;
            end
            if(_zz_8) begin
              buffer_array_2_data_0_1 <= out_MatZ_Bundle_wire_0_1_data;
            end
          end
          if(out_MatZ_Bundle_wire_1_0_Final) begin
            if(_zz_6) begin
              buffer_array_0_data_1_0 <= out_MatZ_Bundle_wire_1_0_data;
            end
            if(_zz_7) begin
              buffer_array_1_data_1_0 <= out_MatZ_Bundle_wire_1_0_data;
            end
            if(_zz_8) begin
              buffer_array_2_data_1_0 <= out_MatZ_Bundle_wire_1_0_data;
            end
          end
          if(out_MatZ_Bundle_wire_1_1_Final) begin
            if(_zz_6) begin
              buffer_array_0_data_1_1 <= out_MatZ_Bundle_wire_1_1_data;
            end
            if(_zz_7) begin
              buffer_array_1_data_1_1 <= out_MatZ_Bundle_wire_1_1_data;
            end
            if(_zz_8) begin
              buffer_array_2_data_1_1 <= out_MatZ_Bundle_wire_1_1_data;
            end
          end
          if(buffer_array_1_Valid) begin
            buffer_array_1_Valid <= 1'b0;
            buffer_array_1_Occupied <= 1'b0;
          end
        end
        if(buffer_array_2_Occupied) begin
          if(out_MatZ_Bundle_wire_0_2_Final) begin
            if(_zz_10) begin
              buffer_array_0_data_0_2 <= out_MatZ_Bundle_wire_0_2_data;
            end
            if(_zz_11) begin
              buffer_array_1_data_0_2 <= out_MatZ_Bundle_wire_0_2_data;
            end
            if(_zz_12) begin
              buffer_array_2_data_0_2 <= out_MatZ_Bundle_wire_0_2_data;
            end
          end
          if(out_MatZ_Bundle_wire_1_2_Final) begin
            if(_zz_10) begin
              buffer_array_0_data_1_2 <= out_MatZ_Bundle_wire_1_2_data;
            end
            if(_zz_11) begin
              buffer_array_1_data_1_2 <= out_MatZ_Bundle_wire_1_2_data;
            end
            if(_zz_12) begin
              buffer_array_2_data_1_2 <= out_MatZ_Bundle_wire_1_2_data;
            end
          end
          if(out_MatZ_Bundle_wire_2_0_Final) begin
            if(_zz_10) begin
              buffer_array_0_data_2_0 <= out_MatZ_Bundle_wire_2_0_data;
            end
            if(_zz_11) begin
              buffer_array_1_data_2_0 <= out_MatZ_Bundle_wire_2_0_data;
            end
            if(_zz_12) begin
              buffer_array_2_data_2_0 <= out_MatZ_Bundle_wire_2_0_data;
            end
          end
          if(out_MatZ_Bundle_wire_2_1_Final) begin
            if(_zz_10) begin
              buffer_array_0_data_2_1 <= out_MatZ_Bundle_wire_2_1_data;
            end
            if(_zz_11) begin
              buffer_array_1_data_2_1 <= out_MatZ_Bundle_wire_2_1_data;
            end
            if(_zz_12) begin
              buffer_array_2_data_2_1 <= out_MatZ_Bundle_wire_2_1_data;
            end
          end
          if(out_MatZ_Bundle_wire_2_2_Final) begin
            if(_zz_10) begin
              buffer_array_0_data_2_2 <= out_MatZ_Bundle_wire_2_2_data;
            end
            if(_zz_11) begin
              buffer_array_1_data_2_2 <= out_MatZ_Bundle_wire_2_2_data;
            end
            if(_zz_12) begin
              buffer_array_2_data_2_2 <= out_MatZ_Bundle_wire_2_2_data;
            end
          end
          if(buffer_array_2_Valid) begin
            buffer_array_2_Valid <= 1'b0;
            buffer_array_2_Occupied <= 1'b0;
          end
        end
      end
    end
  end


endmodule
